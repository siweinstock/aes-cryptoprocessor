module sbox (i, o);
    input [7:0] i;
    output [7:0] o;

    reg [7:0] o;

    always @(i) begin
        case (i)
            8'h00: o = 8'h63;
            8'h01: o = 8'h7c;
            8'h02: o = 8'h77;
            8'h03: o = 8'h7b;
            8'h04: o = 8'hf2;
            8'h05: o = 8'h6b;
            8'h06: o = 8'h6f;
            8'h07: o = 8'hc5;
            8'h08: o = 8'h30;
            8'h09: o = 8'h1;
            8'h0A: o = 8'h67;
            8'h0B: o = 8'h2b;
            8'h0C: o = 8'hfe;
            8'h0D: o = 8'hd7;
            8'h0E: o = 8'hab;
            8'h0F: o = 8'h76;
            8'h10: o = 8'hca;
            8'h11: o = 8'h82;
            8'h12: o = 8'hc9;
            8'h13: o = 8'h7d;
            8'h14: o = 8'hfa;
            8'h15: o = 8'h59;
            8'h16: o = 8'h47;
            8'h17: o = 8'hf0;
            8'h18: o = 8'had;
            8'h19: o = 8'hd4;
            8'h1A: o = 8'ha2;
            8'h1B: o = 8'haf;
            8'h1C: o = 8'h9c;
            8'h1D: o = 8'ha4;
            8'h1E: o = 8'h72;
            8'h1F: o = 8'hc0;
            8'h20: o = 8'hb7;
            8'h21: o = 8'hfd;
            8'h22: o = 8'h93;
            8'h23: o = 8'h26;
            8'h24: o = 8'h36;
            8'h25: o = 8'h3f;
            8'h26: o = 8'hf7;
            8'h27: o = 8'hcc;
            8'h28: o = 8'h34;
            8'h29: o = 8'ha5;
            8'h2A: o = 8'he5;
            8'h2B: o = 8'hf1;
            8'h2C: o = 8'h71;
            8'h2D: o = 8'hd8;
            8'h2E: o = 8'h31;
            8'h2F: o = 8'h15;
            8'h30: o = 8'h4;
            8'h31: o = 8'hc7;
            8'h32: o = 8'h23;
            8'h33: o = 8'hc3;
            8'h34: o = 8'h18;
            8'h35: o = 8'h96;
            8'h36: o = 8'h5;
            8'h37: o = 8'h9a;
            8'h38: o = 8'h7;
            8'h39: o = 8'h12;
            8'h3A: o = 8'h80;
            8'h3B: o = 8'he2;
            8'h3C: o = 8'heb;
            8'h3D: o = 8'h27;
            8'h3E: o = 8'hb2;
            8'h3F: o = 8'h75;
            8'h40: o = 8'h9;
            8'h41: o = 8'h83;
            8'h42: o = 8'h2c;
            8'h43: o = 8'h1a;
            8'h44: o = 8'h1b;
            8'h45: o = 8'h6e;
            8'h46: o = 8'h5a;
            8'h47: o = 8'ha0;
            8'h48: o = 8'h52;
            8'h49: o = 8'h3b;
            8'h4A: o = 8'hd6;
            8'h4B: o = 8'hb3;
            8'h4C: o = 8'h29;
            8'h4D: o = 8'he3;
            8'h4E: o = 8'h2f;
            8'h4F: o = 8'h84;
            8'h50: o = 8'h53;
            8'h51: o = 8'hd1;
            8'h52: o = 8'h0;
            8'h53: o = 8'hed;
            8'h54: o = 8'h20;
            8'h55: o = 8'hfc;
            8'h56: o = 8'hb1;
            8'h57: o = 8'h5b;
            8'h58: o = 8'h6a;
            8'h59: o = 8'hcb;
            8'h5A: o = 8'hbe;
            8'h5B: o = 8'h39;
            8'h5C: o = 8'h4a;
            8'h5D: o = 8'h4c;
            8'h5E: o = 8'h58;
            8'h5F: o = 8'hcf;
            8'h60: o = 8'hd0;
            8'h61: o = 8'hef;
            8'h62: o = 8'haa;
            8'h63: o = 8'hfb;
            8'h64: o = 8'h43;
            8'h65: o = 8'h4d;
            8'h66: o = 8'h33;
            8'h67: o = 8'h85;
            8'h68: o = 8'h45;
            8'h69: o = 8'hf9;
            8'h6A: o = 8'h2;
            8'h6B: o = 8'h7f;
            8'h6C: o = 8'h50;
            8'h6D: o = 8'h3c;
            8'h6E: o = 8'h9f;
            8'h6F: o = 8'ha8;
            8'h70: o = 8'h51;
            8'h71: o = 8'ha3;
            8'h72: o = 8'h40;
            8'h73: o = 8'h8f;
            8'h74: o = 8'h92;
            8'h75: o = 8'h9d;
            8'h76: o = 8'h38;
            8'h77: o = 8'hf5;
            8'h78: o = 8'hbc;
            8'h79: o = 8'hb6;
            8'h7A: o = 8'hda;
            8'h7B: o = 8'h21;
            8'h7C: o = 8'h10;
            8'h7D: o = 8'hff;
            8'h7E: o = 8'hf3;
            8'h7F: o = 8'hd2;
            8'h80: o = 8'hcd;
            8'h81: o = 8'h0c;
            8'h82: o = 8'h13;
            8'h83: o = 8'hec;
            8'h84: o = 8'h5f;
            8'h85: o = 8'h97;
            8'h86: o = 8'h44;
            8'h87: o = 8'h17;
            8'h88: o = 8'hc4;
            8'h89: o = 8'ha7;
            8'h8A: o = 8'h7e;
            8'h8B: o = 8'h3d;
            8'h8C: o = 8'h64;
            8'h8D: o = 8'h5d;
            8'h8E: o = 8'h19;
            8'h8F: o = 8'h73;
            8'h90: o = 8'h60;
            8'h91: o = 8'h81;
            8'h92: o = 8'h4f;
            8'h93: o = 8'hdc;
            8'h94: o = 8'h22;
            8'h95: o = 8'h2a;
            8'h96: o = 8'h90;
            8'h97: o = 8'h88;
            8'h98: o = 8'h46;
            8'h99: o = 8'hee;
            8'h9A: o = 8'hb8;
            8'h9B: o = 8'h14;
            8'h9C: o = 8'hde;
            8'h9D: o = 8'h5e;
            8'h9E: o = 8'h0b;
            8'h9F: o = 8'hdb;
            8'hA0: o = 8'he0;
            8'hA1: o = 8'h32;
            8'hA2: o = 8'h3a;
            8'hA3: o = 8'h0a;
            8'hA4: o = 8'h49;
            8'hA5: o = 8'h6;
            8'hA6: o = 8'h24;
            8'hA7: o = 8'h5c;
            8'hA8: o = 8'hc2;
            8'hA9: o = 8'hd3;
            8'hAA: o = 8'hac;
            8'hAB: o = 8'h62;
            8'hAC: o = 8'h91;
            8'hAD: o = 8'h95;
            8'hAE: o = 8'he4;
            8'hAF: o = 8'h79;
            8'hB0: o = 8'he7;
            8'hB1: o = 8'hc8;
            8'hB2: o = 8'h37;
            8'hB3: o = 8'h6d;
            8'hB4: o = 8'h8d;
            8'hB5: o = 8'hd5;
            8'hB6: o = 8'h4e;
            8'hB7: o = 8'ha9;
            8'hB8: o = 8'h6c;
            8'hB9: o = 8'h56;
            8'hBA: o = 8'hf4;
            8'hBB: o = 8'hea;
            8'hBC: o = 8'h65;
            8'hBD: o = 8'h7a;
            8'hBE: o = 8'hae;
            8'hBF: o = 8'h8;
            8'hC0: o = 8'hba;
            8'hC1: o = 8'h78;
            8'hC2: o = 8'h25;
            8'hC3: o = 8'h2e;
            8'hC4: o = 8'h1c;
            8'hC5: o = 8'ha6;
            8'hC6: o = 8'hb4;
            8'hC7: o = 8'hc6;
            8'hC8: o = 8'he8;
            8'hC9: o = 8'hdd;
            8'hCA: o = 8'h74;
            8'hCB: o = 8'h1f;
            8'hCC: o = 8'h4b;
            8'hCD: o = 8'hbd;
            8'hCE: o = 8'h8b;
            8'hCF: o = 8'h8a;
            8'hD0: o = 8'h70;
            8'hD1: o = 8'h3e;
            8'hD2: o = 8'hb5;
            8'hD3: o = 8'h66;
            8'hD4: o = 8'h48;
            8'hD5: o = 8'h3;
            8'hD6: o = 8'hf6;
            8'hD7: o = 8'h0e;
            8'hD8: o = 8'h61;
            8'hD9: o = 8'h35;
            8'hDA: o = 8'h57;
            8'hDB: o = 8'hb9;
            8'hDC: o = 8'h86;
            8'hDD: o = 8'hc1;
            8'hDE: o = 8'h1d;
            8'hDF: o = 8'h9e;
            8'hE0: o = 8'he1;
            8'hE1: o = 8'hf8;
            8'hE2: o = 8'h98;
            8'hE3: o = 8'h11;
            8'hE4: o = 8'h69;
            8'hE5: o = 8'hd9;
            8'hE6: o = 8'h8e;
            8'hE7: o = 8'h94;
            8'hE8: o = 8'h9b;
            8'hE9: o = 8'h1e;
            8'hEA: o = 8'h87;
            8'hEB: o = 8'he9;
            8'hEC: o = 8'hce;
            8'hED: o = 8'h55;
            8'hEE: o = 8'h28;
            8'hEF: o = 8'hdf;
            8'hF0: o = 8'h8c;
            8'hF1: o = 8'ha1;
            8'hF2: o = 8'h89;
            8'hF3: o = 8'h0d;
            8'hF4: o = 8'hbf;
            8'hF5: o = 8'he6;
            8'hF6: o = 8'h42;
            8'hF7: o = 8'h68;
            8'hF8: o = 8'h41;
            8'hF9: o = 8'h99;
            8'hFA: o = 8'h2d;
            8'hFB: o = 8'h0f;
            8'hFC: o = 8'hb0;
            8'hFD: o = 8'h54;
            8'hFE: o = 8'hbb;
            8'hFF: o = 8'h16;
            default: o = 8'h00;
        endcase
    end

endmodule